library IEEE;
use IEEE.std_logic_1164.all; --  libreria IEEE con definizione tipi standard logic
use WORK.constants.all; -- libreria WORK user-defined

--entity MUX21 is
--        generic( 
--	Port (	A:	In	std_logic;
--		B:	In	std_logic;
--		S:	In	std_logic;
--		Y:	Out	std_logic);
--end MUX21;


entity MUX21_GENERIC IS
	Generic (NBIT: integer:= numBit;
		 DELAY_MUX: Time:= tp_mux);
	Port (	A:	In	std_logic_vector(NBIT-1 downto 0) ;
		B:	In	std_logic_vector(NBIT-1 downto 0);
		SEL:	In	std_logic;
		Y:	Out	std_logic_vector(NBIT-1 downto 0));
	end MUX21_GENERIC;




architecture BEHAVIORAL_5 of MUX21_GENERIC is
begin
	process(A,B,SEL)
	begin
		if (SEL='1') then
			--Y <= A after DELAY_MUX;
                        Y <= A;
		else
			--Y <= B after DELAY_MUX;
                        Y <= B;
		end if;

	end process;

end BEHAVIORAL_5;



architecture STRUCTURAL of MUX21_GENERIC is

	signal Y1: std_logic_vector(NBIT-1 downto 0);
	signal Y2: std_logic_vector(NBIT-1 downto 0);
	signal SB: std_logic;

	component ND2
	Port (	A:	In	std_logic;
		B:	In	std_logic;
		Y:	Out	std_logic);
	end component;
	
	component IV
	Port (	A:	In	std_logic;
		Y:	Out	std_logic);
	end component;

begin


UIV : IV
	Port Map ( SEL, SB);

UND1 : for i in 0 to NBIT-1 generate
       begin 
	    UND1_i : ND2
	    Port Map ( A(i), SEL, Y1(i));
	end generate;

UND2 : for i in 0 to NBIT-1 generate
       begin
            UND2_i : ND2
            Port Map ( B(i), SB, Y2(i));
       end generate;

UND3 : for i in 0 to NBIT-1 generate
       begin
            UND3_i : ND2
	    Port Map ( Y1(i), Y2(i), Y(i));
        end generate;

end STRUCTURAL;




configuration CFG_MUX21_GEN_BEHAVIORAL of MUX21_GENERIC is
	for BEHAVIORAL_5
	end for;
end CFG_MUX21_GEN_BEHAVIORAL;

configuration CFG_MUX21_GEN_STRUCTURAL of MUX21_GENERIC is
	for STRUCTURAL
		for all : IV
			use configuration WORK.CFG_IV_BEHAVIORAL;
		end for;
		for all : ND2
			use configuration WORK.CFG_ND2_ARCH2;
		end for;
	end for;
end CFG_MUX21_GEN_STRUCTURAL;
